module register_file (
  //parameters
) (
  //ports
);
  
endmodule